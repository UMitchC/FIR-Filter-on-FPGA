-- usb.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity usb is
	port (
		address    : in    std_logic_vector(1 downto 0)  := (others => '0'); --   avalon_usb_slave.address
		chipselect : in    std_logic                     := '0';             --                   .chipselect
		read       : in    std_logic                     := '0';             --                   .read
		write      : in    std_logic                     := '0';             --                   .write
		writedata  : in    std_logic_vector(15 downto 0) := (others => '0'); --                   .writedata
		readdata   : out   std_logic_vector(15 downto 0);                    --                   .readdata
		clk        : in    std_logic                     := '0';             --                clk.clk
		OTG_INT1   : in    std_logic                     := '0';             -- external_interface.INT1
		OTG_DATA   : inout std_logic_vector(15 downto 0) := (others => '0'); --                   .DATA
		OTG_RST_N  : out   std_logic;                                        --                   .RST_N
		OTG_ADDR   : out   std_logic_vector(1 downto 0);                     --                   .ADDR
		OTG_CS_N   : out   std_logic;                                        --                   .CS_N
		OTG_RD_N   : out   std_logic;                                        --                   .RD_N
		OTG_WR_N   : out   std_logic;                                        --                   .WR_N
		OTG_INT0   : in    std_logic                     := '0';             --                   .INT0
		irq        : out   std_logic;                                        --          interrupt.irq
		reset      : in    std_logic                     := '0'              --              reset.reset
	);
end entity usb;

architecture rtl of usb is
	component usb_usb_0 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset      : in    std_logic                     := 'X';             -- reset
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect : in    std_logic                     := 'X';             -- chipselect
			read       : in    std_logic                     := 'X';             -- read
			write      : in    std_logic                     := 'X';             -- write
			writedata  : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out   std_logic_vector(15 downto 0);                    -- readdata
			irq        : out   std_logic;                                        -- irq
			OTG_INT1   : in    std_logic                     := 'X';             -- export
			OTG_DATA   : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			OTG_RST_N  : out   std_logic;                                        -- export
			OTG_ADDR   : out   std_logic_vector(1 downto 0);                     -- export
			OTG_CS_N   : out   std_logic;                                        -- export
			OTG_RD_N   : out   std_logic;                                        -- export
			OTG_WR_N   : out   std_logic;                                        -- export
			OTG_INT0   : in    std_logic                     := 'X'              -- export
		);
	end component usb_usb_0;

begin

	usb_0 : component usb_usb_0
		port map (
			clk        => clk,        --                clk.clk
			reset      => reset,      --              reset.reset
			address    => address,    --   avalon_usb_slave.address
			chipselect => chipselect, --                   .chipselect
			read       => read,       --                   .read
			write      => write,      --                   .write
			writedata  => writedata,  --                   .writedata
			readdata   => readdata,   --                   .readdata
			irq        => irq,        --          interrupt.irq
			OTG_INT1   => OTG_INT1,   -- external_interface.export
			OTG_DATA   => OTG_DATA,   --                   .export
			OTG_RST_N  => OTG_RST_N,  --                   .export
			OTG_ADDR   => OTG_ADDR,   --                   .export
			OTG_CS_N   => OTG_CS_N,   --                   .export
			OTG_RD_N   => OTG_RD_N,   --                   .export
			OTG_WR_N   => OTG_WR_N,   --                   .export
			OTG_INT0   => OTG_INT0    --                   .export
		);

end architecture rtl; -- of usb
