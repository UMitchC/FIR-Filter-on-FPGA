module fftpga (              
	input                     sys_clk,
	input                     sys_rst,
	//////////////
	//audio part//
	//////////////
	//WM978 interface
	input                     aud_bclk,   //bit clk
	input                     aud_lrc,    //synchronize signal
	input                     aud_adcdat, //audio_input
	input                     key0,
	output                    aud_mclk,   //main clk signal for WM8978,generated by pll ip core
	output                    aud_dacdat,  //audio output
	//control interface
	output                    aud_scl,    //WM8978 audio IIC clock signal
	inout                     aud_sda    //WM8978 audio IIC data signal
);

//parameter define


//reg define

//wire define
wire    [15:0]      adc_data;   //audio data sampled by FPGA
wire    [33:0]      fir_data;   //audio output form the fir filter
wire                rx_done;    //an output from the audio interface
//signals connecting the fft module and the lcd_top module
wire    [15:0]      audio_data_out; //the data going to the wm8978 input port

//************************************************************************************
//                 main code
//************************************************************************************
//assign audio_data_out = key0?adc_data:fir_data[33:18]; //if press the button key0 then output is filtered data
//the audio part
//the pll module is just to generate a 12MHz signal and to be the main clock signal of the chip
pll_clk u_pll_clk(
    .areset             (~sys_rst  ),   
    .inclk0             (sys_clk   ),   
    .c0                 (aud_mclk  )    //the output to be the clock of the chip
);

//WM8978 control
wm8978_ctrl u_wm8978_ctrl(
    .clk                (sys_clk    ),  
    .rst_n              (sys_rst    ),  

    .aud_bclk           (aud_bclk   ),  //clk signal coming from the chip, control the data transmission
    .aud_lrc            (aud_lrc    ),  //synchronization signal
    .aud_adcdat         (aud_adcdat ),  //data transmission
    .aud_dacdat         (aud_dacdat ),  
    
    .aud_scl            (aud_scl    ),  //scl signal of IIC
    .aud_sda            (aud_sda    ),  //SDA signal of IIC
    
    .adc_data           (adc_data   ),  
    .dac_data           (audio_data_out   ),  /////////need to be changed to fir_data//////////////////////////
    .rx_done            (rx_done),             
    .tx_done            ()              
);



//fir filter module, get data from the receiver and do filtering
fir_filter_mat u_fir_filter_mat(
	 .clk            (aud_bclk),
	 .reset          (sys_rst),
	 //audio input 
	 .clk_enable     (rx_done),
	 .filter_in       (adc_data),
	 //output signals
	 .filter_out      (fir_data),

);


select u_select(
	//input signal
	.key0							(key0),
	.adc_data				   (adc_data),	
	.fir_data               (fir_data[33:18]),
	//output signal
	.audio_data_out			(audio_data_out)
);
endmodule
